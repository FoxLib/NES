// Модуль видеоадаптера

module ppu(

    // 25 мегагерц
    input   wire        clock,      // Входящий 25 Мгц
    output  reg         clock_ppu,  // Тактовый сигнал PPU
    output  wire        clock_cpu,  // Chip Enable для CPU

    // Подключение к видеопамяти
    output reg [10:0]   cursor,
    output reg [12:0]   cursor_chr,
    output reg [ 7:0]   cursor_oam,
    input  wire [7:0]   data,
    input  wire [7:0]   data_chr,
    input  wire [7:0]   data_oam,

    // Выходные данные
    output  reg  [3:0]  r,
    output  reg  [3:0]  g,
    output  reg  [3:0]  b,
    output  wire        hs,
    output  wire        vs
);

// Берется лишь 1 такт из 25 Мгц диапазона для CPU
assign clock_cpu = (cpu_cnt == 2'b01) && clock_ppu && ~clock;

//======================================================================
//  Тактовый генератор
//           ___     ___     ___     ___     ___     ___     ___     ___
// CLK25 ___|///|___|///|___|///|___|///|___|///|___|///|___|///|___|///
//           _______         _______         _______         _______
// PPU   ___|///////|_______|///////|_______|///////|_______|///////|___
// cnt =  0 | 1             | 2             | 0             | 1
//          ^ ppu clock
//               ___                                             ___
// CPU   _______|///|___________________________________________|///|___
//                   ^ cpu clock
//
//======================================================================

initial begin

    clock_ppu = 0;

    // Unchained
    // BG: 0F 0C 1C 30 | 0F 0C 28 38 | 0F 0C 1C 2C | 0F 0C 0F 1C
    // SP: 00 06 16 26 | 0F 0F 18 28 | 0F 01 00 30 | 0F 30 38 16

    // Mario
    // BG: 22 29 1A 0F | 0F 36 17 0F | 0F 30 21 0F | 0F 27 17 0F
    // SP: 00 16 27 18 | 0F 1A 30 27 | 0F 16 30 27 | 0F 0F 36 17

    /* 0 */  Palette_BG[0]  = 6'h22;   Palette_SP[0]  = 6'h00;
    /* 1 */  Palette_BG[1]  = 6'h29;   Palette_SP[1]  = 6'h16;
    /* 2 */  Palette_BG[2]  = 6'h1A;   Palette_SP[2]  = 6'h27;
    /* 3 */  Palette_BG[3]  = 6'h0F;   Palette_SP[3]  = 6'h18;

    /* 4 */
    /* 5 */  Palette_BG[5]  = 6'h36;   Palette_SP[5]  = 6'h1A;
    /* 6 */  Palette_BG[6]  = 6'h17;   Palette_SP[6]  = 6'h30;
    /* 7 */  Palette_BG[7]  = 6'h0F;   Palette_SP[7]  = 6'h27;

    /* 8 */
    /* 9 */  Palette_BG[9]  = 6'h30;   Palette_SP[9]  = 6'h16;
    /* 10 */ Palette_BG[10] = 6'h21;   Palette_SP[10] = 6'h30;
    /* 11 */ Palette_BG[11] = 6'h0F;   Palette_SP[11] = 6'h27;

    /* 12 */
    /* 13 */ Palette_BG[13] = 6'h27;   Palette_SP[13] = 6'h0F;
    /* 14 */ Palette_BG[14] = 6'h17;   Palette_SP[14] = 6'h36;
    /* 15 */ Palette_BG[15] = 6'h0F;   Palette_SP[15] = 6'h17;

    // Курсоры
    cursor     = 0;
    cursor_chr = 0;
    cursor_oam = 0;

    // Спрайты (для теста)
    sprites_temp[0] = 32'h00_00_00_00;
    sprites_temp[1] = 32'h00_00_00_00;
    sprites_temp[2] = 32'h00_00_00_00;
    sprites_temp[3] = 32'h00_00_00_00;
    sprites_temp[4] = 32'h00_00_00_00;
    sprites_temp[5] = 32'h00_00_00_00;
    sprites_temp[6] = 32'h00_00_00_00;
    sprites_temp[7] = 32'h00_00_00_00;

end

// Тайминги для горизонтальной развертки (640)
parameter horiz_visible = 640;
parameter horiz_back    = 48;
parameter horiz_sync    = 96;
parameter horiz_front   = 16;
parameter horiz_whole   = 800;

// Тайминги для вертикальной развертки (480)
//                              // 400  480
parameter vert_visible = 480;   // 400  480
parameter vert_back    = 33;    // 35   33
parameter vert_sync    = 2;     // 2    2
parameter vert_front   = 10;    // 12   10
parameter vert_whole   = 525;   // 449  525

// Начало и конец области рисования
parameter start_x      = 64 - 16;
parameter end_x        = start_x + 512 + 16;

// 640 (видимая область) + 48 (задний порожек) + 96 (синхронизация) + 16 (передний порожек)
assign hs = x >= (640 + horiz_front) && x < (640 + horiz_front + horiz_sync);
assign vs = y >= (480 + vert_front)  && y < (480 + vert_front  + vert_sync);

// Текущее положение луча на экране
reg  [9:0] x = 1'b0;
reg  [9:0] y = 1'b0;

// Делитель CPU [0,1,2]
reg  [1:0] cpu_cnt   = 2'b00;

// ---------------------------------------------------------------------
//  Регистры контроля
// ---------------------------------------------------------------------

                  ///  7 65 43 2 10
reg [7:0]  CTRL0  = 8'b0_00_10_0_00;

/*
7   Формирование запроса прерывания NMI при кадровом синхроимпульсе
    (0 - запрещено; 1 - разрешено)

6   (Не используется, должен быть 0)
5   Размер спрайтов (0 - 8x8; 1 - 8x16)
4   Выбор знакогенератора фона (0/1)
3   Выбор знакогенератора спрайтов (0/1)
2   Выбор режима инкремента адреса при обращении к видеопамяти
    (0 – увеличение на единицу «горизонтальная запись»;
     1 - увеличение на 32 «вертикальная запись»)

1,0 Адрес активной экранной страницы
    (00 – $2000; 01 – $2400; 10 – $2800; 11 - $2C00)
*/

//                     76543210
reg [7:0]  CTRL1  = 8'b00011000;

/* 7-5     Яркость экрана/интенсивность цвета в RGB (в Денди не используется)
    4      0 – Спрайты не отображаются; 1 – Спрайты отображаются
    3      0 – Фон не отображается; 1 – Фон отображается
    2      0 – Спрайты невидны в крайнем левом столбце; 1- Все спрайты видны
    1      0 – Рисунок фона невиден в крайнем левом столбце; 1 - Весь фон виден
    0      Тип дисплея: Color/Monochrome (в Денди не используется) */

// ---------------------------------------------------------------------
// Регистры для отрисовки изображения на экране
// ---------------------------------------------------------------------

reg  [1:0]  NTA     = 2'b00;
wire        NTBank  = NTA[0] ^ NTA[1] ^ X[8] ^ RegH ^ RegV;

// Текущее положение луча
reg  [8:0]  PPUX    = 9'h0;  /* 0..340 */
reg  [8:0]  PPUY    = 9'h0;  /* 0..261 */

// Калибровочные скроллинги
reg         RegH    = 0; // Смена страницы по X
reg         RegV    = 0; // Смена страницы по Y
reg  [4:0]  RegHT   = 0; // Грубый горизонтальный
reg  [4:0]  RegVT   = 0; // Грубый вертикальный
reg  [3:0]  RegFH   = 0; // Точный горизонтальный
reg  [3:0]  RegFV   = 0; // Точный вертикальный

// Положение пера для рисования на холсте 256x240
wire [8:0] X = PPUX[8:0] + {RegHT[4:0], RegFH[2:0]} - 8;
wire [8:0] Y = PPUY[8:0] + {RegVT[4:0], RegFV[2:0]};

/* Цветовые атрибуты фона */
reg  [7:0]  chrl;       /* Нижние  8 бит цвета */
reg  [7:0]  chrh;       /* Старшие 8 бит цвета */
reg  [7:0]  hiclr;      /* 3=[7:6] 2=[5:4] 1=[3:2] 0=[1:0] */
reg  [1:0]  colorpad;   /* Атрибуты */
reg  [15:0] colormap;   /* Цвета битов */

/* Палитры в регистрах PPU */
reg  [ 5:0] Palette_BG[16];  /* Палитра фона */
reg  [ 5:0] Palette_SP[16];  /* Палитра спрайтов */
reg  [5:0]  color;           /* Текущий цвет из глобальной палитры */
reg  [15:0] rgb;             /* Реальный VGA-цвет */

/* Спрайты */
// ---------------------------------------------------------------------

// Временное хранилище для спрайтов, которые собираются из памяти OAM
// при сканировании очередной линии

/*
 31:24 Y        | CHR-HI
 23:16 Attrs
 15:8  SpriteID | CHR-LOW
  7:0  X
*/

reg  [31:0] sprites_temp [8]; // Временно
reg  [31:0] sprites      [8]; // Постоянно

// Каждый бит в `sp_live` говорит о том, будет ли использован sprites[n]
// для рисования, или нет. Это нужно чтобы не отображать на экране не
// используемые спрайты

reg  [ 7:0] sp_live_temp = 8'h00; // Временное хранилище
reg  [ 7:0] sp_live      = 8'h00; // Не изменяется на следующей линии

// Важный параметр. Zero-спрайт. Если такой спрайт находится на линии,
// это значит, что будет возведен особый флаг Sprite0Hit, который будет
// сигнализировать о достижении лучом нулевого спрайта. Обрабатывается
// отдельно
reg         sp_zero_temp = 1'b0;
reg         sp_zero      = 1'b0;

// Счетчик спрайтов. Если он достиг >7, то более не добавляется в sp_hits
// и также не добавляется в sprites_temp при вычислении
reg  [ 3:0] sp_counter = 0;
reg         sp_hit     = 0; // Если sp_hit=1 то значит, что спрайт ПОПАЛ в область видимости
reg  [ 2:0] sp_icon_id = 7; // Иконка, у которой необходимо получить атрибуты из CHR-ROM

// Идентификатор иконки у спрайта (какую иконку он использует)
wire [7:0]  sp_icon    = sprites_temp[ sp_icon_id ][ 15:8 ];

// Отражения спрайта
wire VMirror = sprites_temp[ sp_icon_id ][ 16 + 7 ]; // Отражение по вертикали?
wire HMirror = sprites_temp[ sp_icon_id ][ 16 + 6 ]; // Отражение по горизонтали?

// Положение внутри спрайта (от 0 до 7/15)
wire [3:0] Ydiff = sprites_temp[ sp_icon_id ][ 27:24 ];

// Реальное положение в зависимости от зеркалирования и размера спрайта
wire [3:0] YVert = VMirror ? ((CTRL0[5] ? 15 : 7) - Ydiff) : Ydiff;

// Зеркалирование по X (если задан параметр)
wire [7:0] FMirr = HMirror ? {data_chr[0], data_chr[1], data_chr[2], data_chr[3], data_chr[4], data_chr[5], data_chr[6], data_chr[7]} : data_chr[7:0];

// ---------------------------------------------------------------------
// Пересчет спрайтов и вычисление конечного цвета
// ---------------------------------------------------------------------

wire [4:0] chain_color[8]; // Вычисления цветов через eval
wire [8:0] sp_x         = PPUX - 16;
wire [7:0] sp_hit_z;    /* Фиксация попадания луча на рисуемый пиксель */
reg  [3:0] bgcolor;     /* Реальный отображаемый цвет фона */
wire [4:0] final_color  = chain_color[7][4:0]; // Последний цвет из спрайтов

/* Текущий рисуемый цвет фона */
wire [3:0] current_bgcolor =
{
    colorpad[            1:0 ], // 2 bit
    colormap[ {X[2:0], 1'b1} ], // 1 bit
    colormap[ {X[2:0], 1'b0} ]  // 1 bit
};

// Вычисление цвета фона
always @* begin

    /* Прозрачный */
    if (current_bgcolor[1:0] == 2'b00)
        bgcolor = 0;

    /* Скрытие левого столбца или всего фона */
    else if ((x < (start_x+32) && CTRL1[1] == 1'b0) || (CTRL1[3] == 1'b0))
        bgcolor = 0;

    /* Реальный цвет */
    else bgcolor = current_bgcolor;

end

// Вычисления спрайтов
//      Упр.   Актуален?   Спрайт      Цвет (вход)     X     Цвет (выход)    Хит лучом
eval S1(CTRL1, sp_live[0], sprites[0], {1'b0,bgcolor}, sp_x, chain_color[0], sp_hit_z[0]);
eval S2(CTRL1, sp_live[1], sprites[1], chain_color[0], sp_x, chain_color[1], sp_hit_z[1]);
eval S3(CTRL1, sp_live[2], sprites[2], chain_color[1], sp_x, chain_color[2], sp_hit_z[2]);
eval S4(CTRL1, sp_live[3], sprites[3], chain_color[2], sp_x, chain_color[3], sp_hit_z[3]);
eval S5(CTRL1, sp_live[4], sprites[4], chain_color[3], sp_x, chain_color[4], sp_hit_z[4]);
eval S6(CTRL1, sp_live[5], sprites[5], chain_color[4], sp_x, chain_color[5], sp_hit_z[5]);
eval S7(CTRL1, sp_live[6], sprites[6], chain_color[5], sp_x, chain_color[6], sp_hit_z[6]);
eval S8(CTRL1, sp_live[7], sprites[7], chain_color[6], sp_x, chain_color[7], sp_hit_z[7]);

/* Решение о том, какой цвет будет выведен */
always @* begin

    /* Если выходит за границы, то цвет будет фоновый в любом случае */
    if (x < (start_x + 16) || x >= (start_x + 512 + 16))
                             color = Palette_BG[ 0 ];
    /* Цвет спрайта */
    else if (final_color[4]) color = Palette_SP[ final_color[3:0] ];
    /* Цвет фона */ else     color = Palette_BG[ final_color[3:0] ];

end

// ---------------------------------------------------------------------
// Базовая частота 25 Мгц
// ---------------------------------------------------------------------

always @(posedge clock) begin

    // -----------------------------------------------------------------
    // Рисование готовых видеоданных на VGA
    // -----------------------------------------------------------------

    if (x < 640 && y < 480) begin

        // Цвет определяется внешним способом
        if (y[0])
            {r, g, b} <= {rgb[4:1], rgb[10:7], rgb[15:12]};
        else
        // Чересстрочная выдача видеоданных
            {r, g, b} <= {1'b0,rgb[4:2],  1'b0,rgb[10:8],  1'b0,rgb[15:13]};

    // Невидимая область
    end else {r, g, b} <= 12'h000;

    // -----------------------------------------------------------------
    // Обработка видимой области
    // A. Чтение символов для видеовыдачи
    // B. Обработка спрайтов (чтение 256 байт из OAM)
    // -----------------------------------------------------------------

    if (x[0]) begin

        // -------------------------------------------------------------
        // Считывание информации спрайтов
        // -------------------------------------------------------------

        // Шаг 1. Защелка спрайтов
        if (PPUX == 0) begin

            // Защелкивание спрайтов
            sp_zero    <= sp_zero_temp;
            sp_live    <= sp_live_temp;
            sprites[0] <= sprites_temp[0];
            sprites[1] <= sprites_temp[1];
            sprites[2] <= sprites_temp[2];
            sprites[3] <= sprites_temp[3];
            sprites[4] <= sprites_temp[4];
            sprites[5] <= sprites_temp[5];
            sprites[6] <= sprites_temp[6];
            sprites[7] <= sprites_temp[7];

            // Инициализация
            sp_live_temp <= 0;
            sp_zero_temp <= 0;

            sp_counter   <= 0;
            cursor_oam   <= 0;

        end

        // Шаг 2. Считывание из OAM
        else if (PPUX >= 8 && PPUX < 9'h108) begin

            case (PPUX[1:0])

            // Проверка на попадание спрайта в диапазон [Y <= PPUY < Y + 8/16]
            // А также НЕ должно быть превышения по количеству одновременных спрайтов
            // на линии (бит sp_counter[3])

            /* +0 Байт Y */
            0: if (~sp_counter[3] && data_oam <= PPUY && PPUY < (data_oam + (CTRL0[5] ? 16 : 8)))
            begin sp_hit <= 1'b1; /* Спрайт виден */

                // Запись Diff для расчета битов по Y
                sprites_temp[ sp_counter[2:0] ][ 31:24 ] <= (PPUY - data_oam);

                // Пишем информацию о том, что спрайт попал в сканлайн
                sp_live_temp[ sp_counter[2:0] ] <= 1'b1;

                // Если это Zero-спрайт, отметить это
                if (cursor_oam == 0) sp_zero_temp <= 1'b1;

            end
            // Спрайт не виден
            else sp_hit <= 1'b0;

            // +1 Загружаем в память иконку спрайта
            2'h1: if (sp_hit) begin sprites_temp[ sp_counter[2:0] ][15:8]  <= data_oam; end

            // +2 Запись атрибутов спрайта
            2'h2: if (sp_hit) begin sprites_temp[ sp_counter[2:0] ][23:16] <= data_oam; end

            // +3 Запись X
            2'h3: if (sp_hit) begin sprites_temp[ sp_counter[2:0] ][7:0] <= data_oam;

                // Переход к следующему спрайту (с учетом что нет overflow)
                if (sp_counter[3] == 0) sp_counter <= sp_counter + 1;

            end
            endcase

            cursor_oam <= cursor_oam + 1;

        end

        // -------------------------------------------------------------
        // Выдача фона и считывание атрибутов спрайтов
        // -------------------------------------------------------------

        // Чтение цветовой маски 8 спрайтов
        if (PPUX >= 9'h108 && PPUX < (9'h108 + 8*4)) begin

            case (PPUX[1:0])

                0: begin sp_icon_id <= PPUX[4:2] - 2; end
                1: begin

                                            //   Банк 0/1    <ID Иконки в банке>     <L/H> Позиция Y
                    if (CTRL0[5]) cursor_chr <= {sp_icon[0], sp_icon[7:1], YVert[3], 1'b0, YVert[2:0]}; // x16
                    else          cursor_chr <= {CTRL0[3],   sp_icon[7:0],           1'b0, YVert[2:0]}; // x8

                end

                // Запись в диапазон, где был +2 ID иконки (теперь там CHR-LOW)
                2: begin sprites_temp[ sp_icon_id ][ 15:8 ]  <= FMirr; cursor_chr[3] <= 1'b1; end

                // Запись в диапазон, где был +0 YDiff (теперь там CHR-HI)
                3: begin sprites_temp[ sp_icon_id ][ 31:24 ] <= FMirr; end

            endcase

        end

        // Чтение знакомест фона
        else case (X[2:0])

            // Прочитаем из памяти символ 8x8
            2'h0: cursor <= {NTBank, Y[7:3], X[7:3]};

            // Начнем чтение CHR (BA=0, CHR=00000000, B=0, Y=000}
            2'h1: begin

                // Чтение младшего бита символа из CHR-ROM
                cursor_chr <= {CTRL0[4], data[7:0], 1'b0, Y[2:0]};

                // Запрос цветовых атрибутов
                cursor     <= {NTBank, 4'b1111, Y[7:5], X[7:5] };

            end

            // Чтение верхней палитры знакогенератора и ATTR
            2'h2: begin

                cursor_chr[3] <= 1'b1; // Установка старшего бита

                hiclr <= data;         // Чтение цветового атрибута
                chrl  <= data_chr;     // Младшие 8 бит цветов из CHR-ROM

            end

            // Прочитаны старшие биты цветов фона
            2'h3: begin chrh  <= data_chr; end

            // Результат
            4'h7: begin

                // Старшие цвета пикселей
                colorpad <= {hiclr[ {Y[4], X[4], 1'b1} ],  // 7|5|3|1
                             hiclr[ {Y[4], X[4], 1'b0} ]}; // 6|4|2|0

                // Нижние цвета пикселей /
                colormap <= {/* BIT 7 */ chrh[0], chrl[0], /* BIT 6 */ chrh[1], chrl[1],
                             /* BIT 5 */ chrh[2], chrl[2], /* BIT 4 */ chrh[3], chrl[3],
                             /* BIT 3 */ chrh[4], chrl[4], /* BIT 2 */ chrh[5], chrl[5],
                             /* BIT 1 */ chrh[6], chrl[6], /* BIT 0 */ chrh[7], chrl[7]};

            end

        endcase

    end

    // -----------------------------------------------------------------
    // Процессинг PPU & CPU
    //  64 = Базовая линия
    // -16 = Отступ для предвычисления символа
    //  +2 = Для коррекции на начало X[2:0] = 0
    // -----------------------------------------------------------------

    // Допустимая зона посередине (341Т) и по высоте (262Т)
    if (x >= (start_x-16+2) && x < ((start_x-16+2) + 341*2) && y < 524) begin

        // Раз в 2Т выполнять такт PPU
        if (x[0]) begin

            // Обработка 1 такта PPU от NES (реальный)
            if (~y[0]) begin

                // Памятка:
                // cpu_cnt = 01 >> Только что отработал такт CPU <<
                // cpu_cnt = 10 Данные из CPU не брать
                // cpu_cnt = 00 Данные из CPU не брать

// !!!!!!!!!!!!!!!! ГРЯЗНЫЙ ХАК -----------------------------------------!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!
CTRL1 <= 8'b000_11_00_0;

                // Формирование разрешений такта на CPU
                cpu_cnt <= (cpu_cnt == 2'b10) ? 0 : cpu_cnt + 1;

            end

            // Сдвиг луча Y при достижении края PPUX на этом сканлайне
            PPUY <= (PPUX == 340 && y[0]) ? PPUY + 1 : PPUY;

            // Луч X сдвигать на каждом (!) сканлайне
            PPUX <= (PPUX == 340) ? 0 : PPUX + 1;

        end
        // Сброс PPU(X|Y) в конце
        else if (y == 523) begin PPUX <= 0; PPUY <= 0; end

        // --------------------
        // Делитель частоты PPU
        // --------------------

        clock_ppu <= x[0] & ~y[0];

    end

    // Полное отключение процессинга (CPU & PPU)
    else begin

        clock_ppu <= 0;
        cpu_cnt   <= 0;

    end

    // Видеокадр
    x <= (x == horiz_whole - 1) ? 1'b0 : (x + 1'b1);
    y <= (x == horiz_whole - 1) ? (y == vert_whole - 1 ? 1'b0 : y + 1'b1) : y;

end

// ---------------------------------------------------------------------
// Преобразования номера цвета палитры в реальный (16 bit)
// ---------------------------------------------------------------------

always @* case (color)

    6'd0:  rgb = 16'h73ae;
	6'd1:  rgb = 16'h88c4;
	6'd2:  rgb = 16'ha800;
	6'd3:  rgb = 16'h9808;
	6'd4:  rgb = 16'h7011;
	6'd5:  rgb = 16'h1015;
	6'd6:  rgb = 16'h0014;
	6'd7:  rgb = 16'h004f;
	6'd8:  rgb = 16'h0168;
	6'd9:  rgb = 16'h0220;
	6'd10: rgb = 16'h0280;
	6'd11: rgb = 16'h11e0;
	6'd12: rgb = 16'h59e3;
	6'd16: rgb = 16'hbdf7;
	6'd17: rgb = 16'heb80;
	6'd18: rgb = 16'he9c4;
	6'd19: rgb = 16'hf010;
	6'd20: rgb = 16'hb817;
	6'd21: rgb = 16'h581c;
	6'd22: rgb = 16'h015b;
	6'd23: rgb = 16'h0a79;
	6'd24: rgb = 16'h0391;
	6'd25: rgb = 16'h04a0;
	6'd26: rgb = 16'h0540;
	6'd27: rgb = 16'h3c80;
	6'd28: rgb = 16'h8c00;
	6'd32: rgb = 16'hffff;
	6'd33: rgb = 16'hfde7;
	6'd34: rgb = 16'hfcab;
	6'd35: rgb = 16'hfc54;
	6'd36: rgb = 16'hfbde;
	6'd37: rgb = 16'hb3bf;
	6'd38: rgb = 16'h63bf;
	6'd39: rgb = 16'h3cdf;
	6'd40: rgb = 16'h3dfe;
	6'd41: rgb = 16'h1690;
	6'd42: rgb = 16'h4ee9;
	6'd43: rgb = 16'h9fcb;
	6'd44: rgb = 16'hdf40;
	6'd48: rgb = 16'hffff;
	6'd49: rgb = 16'hff35;
	6'd50: rgb = 16'hfeb8;
	6'd51: rgb = 16'hfe5a;
	6'd52: rgb = 16'hfe3f;
	6'd53: rgb = 16'hde3f;
	6'd54: rgb = 16'hb5ff;
	6'd55: rgb = 16'haedf;
	6'd56: rgb = 16'ha73f;
	6'd57: rgb = 16'ha7fc;
	6'd58: rgb = 16'hbf95;
	6'd59: rgb = 16'hcff6;
	6'd60: rgb = 16'hf7f3;
	default: rgb = 1'b0;

endcase

endmodule
